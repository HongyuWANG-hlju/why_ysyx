`include "defines.v"

module m_stage(
    
);
    
endmodule